module f6();
endmodule
module f1_core1 ();

endmodule
module f1_test();
    endmodule


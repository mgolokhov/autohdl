module f1 ();
endmodule

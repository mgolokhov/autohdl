module f5();
endmodule

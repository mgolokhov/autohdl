module inst3 (input a, input b); endmodule

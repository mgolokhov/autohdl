module f2_dsn1_uncopied();
endmodule

module f1_dsn1 ();

f1_core2 f1_core2_inst();

endmodule

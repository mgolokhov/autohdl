//**********������ ��������� �������������� ������ �������� � ���������*****************************//
//����������: ������ ��������� �������������� ������ �������� � ��������� ��������������� ��� ���������� ������ � �������
//��������� ���� resolver_kalman. ��������! ���� ����������� �� ��������. ���� ����� ������� ����� 2048 ������ �������� �� �����������.
//�����:
//rst	    - ����������� �����
//clk	    - �������� ���������		  
//cA       - ���� �� ������ A
//cB       - ���� �� ������ B
//cC       - ���� �� ������ C (����-�����)
//
//������:
//phi       - ���������, �������� 32 ���. ���������� �������������� ���/��� = pi/2^15
//omega     - ��������, �������� 31 ���.
//to		- �������� ������� ����� ����� �������� � ������(30 ���, �����������)
//phi_rdy   - ���� ���������� ���������
//omega_rdy - ���� ���������� ��������
//sync_rst  - c��������� ����� ����
//																
//������������ ��������� � �������� ���������� 1 ���� ��� ��������� (20 �� ��� clk 50 ���)
//������������ ��������� � �������� ���������� 32 ����� ��� �������� (640 �� ��� clk 50 ���)
//
//�����: ������� �.�.
//		 ������� "������� ����������" �����(��), 2009 �.
//**************************************************************************************************//
module quad_sensor_core(rst,clk,cA,cB,cC,phi,omega,phi_rdy,omega_rdy,sync_rst,to,out,acc_level);
	input  rst;  			//����������� �����
	input  clk;  			//�������� ���������
	input  cA;				//���� �� ������ A
	input  cB;				//���� �� ������ B
	input  cC;				//���� �� ������ C (���� �����)
	output reg[31:0]phi;	//��������� �� ������� pi[���] = 2^15. (32 ����, ��������)
	output reg[30:0]omega;	//�������� �� �������  (31 ���, ��������)
	output reg[29:0]to;		//�������� ������� ����� ����� �������� � ������(30 ���, �����������)	  
	input  [15:0]acc_level;
	output reg[15:0]out;	
	
	output reg phi_rdy;		//�������� ��������� ����������
	output reg omega_rdy;	//�������� �������� ����������			 					 
	output reg sync_rst;	//���������� ����� ���� �� ����� ������� 0 �����
	
parameter ZeroPHI=32'h0;	
parameter ZeroSpeedN = 24;  //����� ���� ���� �������� �������� �� �������������. �.� �� ���������, ��� ���� �� ���� ����� � ������� 2^25 ������, �� �������� ����� 0

reg p_A; 	//���������� �������� ������ A
reg p_B;	//���������� �������� ������ B
reg p_C;	//���������� �������� ������ C	 	 
reg dir;	//����������� 1 - �������������, 0 - �������������
reg [30:0]omegaTimer; //������ ��� ������� �������� ������� ����������
reg WasOverflow;		 
 		 

reg  start;
reg  [29:0]t;
wire [29:0]spd;		  

reg  tmp_dir;	//����������� �� ������ ������ ���������� ��������

reg [30:0]nomega;

always @(*)
	if(tmp_dir)
		nomega<={tmp_dir,-spd};
	else 
		nomega<={tmp_dir,spd};	

wire [31:0]domega;
wire [30:0]abs_domega;

assign domega = {nomega[30],nomega}-{omega[30],omega};
assign abs_domega = domega[31] ? - domega : domega;

wire rdy;

parameter NO_SPEED_LIMIT = 1;  //���� 1, �� ��� ����������� ��������

cordic_inv_t_core inv_t (.rst(rst),
						 .clk(clk),
						 .start(start),
						 .t(t),
						 .spd(spd),
						 .rdy(rdy)
);

reg ch_on_boot;			   

reg chA; 	//�������� ������ A
reg chB;	//�������� ������ B
reg chC;	//�������� ������ C	 	 	   




always @(posedge rst or posedge clk)
	if (rst)
		begin
			chA <= 0;
			chB <= 0;
			chC <= 0;
		end	else
		begin
			chA <= cA;
			chB <= cB;
			chC <= cC;
		end	

always @(posedge rst or posedge clk)
	if(rst)
		begin
			ch_on_boot<=1'b1;
			p_A<=1'b0;
			p_B<=1'b0;
			p_C<=1'b0;						
			omega<=16'd0;	 
			phi<=32'd0;	
			phi_rdy<=1'b0;
			start<=1'b0;
			omega_rdy<=1'b0;
			omegaTimer<=31'd1; //������ ������ � 1, �.�. �� ���� ����� �� ��� �� ����������, � �� ��������� ��� ������� 1 ����
			dir<=1'b0;
			WasOverflow<=1'b0;
			t<=30'd0;	  
			sync_rst<=1'b0;		
			to <=0;
			tmp_dir <= 0;	 
			out<=0;
		end	else
		begin	 
			if (ch_on_boot)
				begin
					ch_on_boot<=1'b0;
					p_A<=chA;
					p_B<=chB;
					p_C<=chC;						
				end			 
			else	
			if ((p_A!=chA)/*||(p_B!=chB)*/)
				begin
					omegaTimer<=31'd1;	//������ ������ � 1, �.�. �� ���� ����� �� ��� �� ����������, � �� ��������� ��� ������� 1 ����
					if (WasOverflow)
						begin																  
							WasOverflow<=1'b0;//������� ���� ������������
							omega<=16'd0;     //���� ���� ���� �� ���� ������������ �������, �� �������� ����� 0
							omega_rdy<=1'b1;  //���������� ����, ���� ��� �������� ���������  
						end	else		 
						begin			 
							if(t[29:12]|(NO_SPEED_LIMIT))	  		  //���� t ����� 2048, �� �������, ��� �������� ��������� �������
								begin 
									start<=1'b1;	  	  //����� �������� ������ �������� ��� 1/omegaTimer*2^30															
									tmp_dir <= dir;
								end	
							to <= omegaTimer[29:0]; //��������� ���������� �������� �������, ���� ��� ��� ������� inv_t_core
                			t<=omegaTimer[29:0]; //��������� ���������� �������� �������, ���� ��� ��� ������� inv_t_core
						end	
				end		
			if ((p_C!=chC))
			begin 		  
				if(chC^dir)
					begin 
						phi<=ZeroPHI;	    //���� ��������� 0 �����, �� ���������� ��������, � ��� ����� ��� ��� ���������
						phi_rdy<=1'b1;	 	//���������� ���� ���������� ���������										   
						sync_rst<=1'b1;
					end
				p_C<=chC;
			end else	
			begin
				sync_rst<=1'b0;
				if (p_A!=chA)			//���� ����� ������ �
					begin	  
						if (chA^chB)
						begin											 
							//************************������������� �����������*******************
							phi[31:14]<=phi[31:14]-1;
							phi_rdy<=1'b1;	 	//���������� ���� ���������� ���������
							dir<=1'b1;			//���������� ��� �����������
							//************************������������� �����������*******************
						end	else
						begin					
							//************************������������� �����������*******************
							phi[31:14]<=phi[31:14]+1;
							phi_rdy<=1'b1;	 	//���������� ���� ���������� ���������
							dir<=1'b0;			//���������� ��� �����������
							//************************������������� �����������*******************
						end		
						p_A<=chA;   //��������� �������� ������ A
					end
				else		
				if (p_B!=chB)
						begin 
							if (chA^chB)
							begin
								//************************������������� �����������*******************
								phi[31:14]<=phi[31:14]+1;
								phi_rdy<=1'b1;	 	//���������� ���� ���������� ���������
								dir<=1'b0;			//���������� ��� �����������
								//************************������������� �����������*******************
							end	else
							begin					
								//************************������������� �����������*******************
								phi[31:14]<=phi[31:14]-1;	
								phi_rdy<=1'b1;	 	//���������� ���� ���������� ���������
								dir<=1'b1;			//���������� ��� �����������
								//************************������������� �����������*******************
							end					
							p_B<=chB;	//��������� �������� ������ B
						end	 else 
						begin			
							to <= {WasOverflow,13'b0,omegaTimer[30:15]}; //��������� ���������� �������� �������, ���� ��� ��� ������� inv_t_core
							phi_rdy<=1'b0;    		//���� ��� ������ ���������� ������ phy_rdy
							if(omegaTimer[ZeroSpeedN])		//���� ������ �������� 30 ���, �� ��������� ������������, ���������� ������ ������� ��� ��� �� ����������
								WasOverflow<=1'b1;
                            else
    							omegaTimer<=omegaTimer+31'd1; //���� �� ���� ������, �� ������������������ ������
						end																					 
			end		
			if (WasOverflow)
				begin 
					omega<=16'd0;     //���� ���� ���� �� ���� ������������ �������, �� �������� ����� 0
					omega_rdy<=1'b1;  //���������� ����, ���� ��� �������� ���������  
				end else
			if (rdy)
				begin					
					if ((abs_domega>{acc_level,4'b0})&(~NO_SPEED_LIMIT))
							out <= out+1;
					else			 
						begin
							omega <= nomega;
							omega_rdy<=1'b1; //���� ������ ����, ����, ��� ������ �������� ����������, �� ������� �� � ������ ����������� � ���������� ���� ���������� �������� ��������
						end
				end else
					if (omega_rdy) omega_rdy<=1'b0; //���� ���� rdy �� ������, � omega_rdy - ���������, �� ������� ���
			if (start) start<=1'b0; //������, ��� ���� ����� ����� ������ ����� �� ��������
		end						 
endmodule

//****************************������ ��������� 19 ���****************************
//
//���-�� ��� ����� ����� - 19 
//�������� ��� - 1
//
//�����:
//a,b - ���������
//������:
//�   - ������������ (�����, �������� 37 ���)						   
//	 
//�����: ������� �.�.
//		 ������� "������� ����������" �����(��), 2009 �.
//********************************************************************************

module mult19(				 
	input  [18:0] a,
	input  [18:0] b,
	output [36:0] c);

wire [18:0]ta_p;    //� ������������ �� -32767 �� 32767
wire [18:0]tb_p;    //b ������������ �� -32767 �� 32767
wire [17:0]ta;      //������ ��������� ta_p           
wire [17:0]tb;	    //������ ��������� tb_p
wire [35:0]mul_res; //��������� ��������� |a|*|b|
wire [35:0]nmul_res;//��������� ��������� |a|*|b| � �������������� ���� ��� ������, ����� a*b<0
wire mul_sign;		//���� ���������			  

assign ta_p		= (a==19'h40000) ? a+1 : a;             
assign tb_p		= (b==19'h40000) ? b+1 : b;
assign ta[17:0] = (ta_p[18]) ? ~ta_p[17:0]+1 : ta_p[17:0];
assign tb[17:0] = (tb_p[18]) ? ~tb_p[17:0]+1 : tb_p[17:0];
assign mul_sign = (ta_p == 19'h0) ? 1'b0 : 
				 ((tb_p == 19'h0) ? 1'b0 : ta_p[18]^tb_p[18]);	
assign c[36]=mul_sign;
assign mul_res=ta*tb;		   
assign nmul_res=-mul_res;
assign c[35:0] = (mul_sign) ? nmul_res[35:0] : mul_res[35:0];

endmodule
module f2 ();


endmodule
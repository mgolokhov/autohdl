module f1 ();
    f2 inst_f2();
endmodule
module top_build_yaml();
endmodule
//***********************************Нечеткий регулятор**************************************************************
//Романов А.М. Кафедра "Проблемы управления" МИРЭА, 2010 г.
//ВАЖНО: x-b+b1, x-b-b1, x-b - для любого a*x[-1:1] окажутся в дипазоне от [-1:1], перед поступлением на умножители, т.к.
//сигмода всегда лежит [0 1]
//а вот x_arg может и не оказаться. Но для s [0 1] вроде как x_arg лежит [-2 2] (надо б еще потестить)
//*******************************************************************************************************************

module fuzzy_PI_cordic
	#(parameter  N=16, 			//Число бит входа и коэффициентов
      parameter  bN=2,           //Число бит целой части b,b1 и s  
      parameter  aN=4           //Число бит целой части a0,a1 
	)	
	(
	input rst,					//Асинхронный сброс
	input clk,					//Тактовый генератор
	input start,				//Строб старта
	input [N-1:0]x,				//Вход x [-1 1]
	input [N-1:0]y,				//Вход y [-1 1]
//(левая функция принадлежноси) 
	input [N-1:0]a0_xl,			//Коэффициент по входу x a0=sqrt(w_x)*sqrt(1-exp(-0.5))/s
	input [N-1:0]a1_xl,			//Коэффициент по входу x a1=sqrt(w_x)*sqrt((1-exp(-0.5))./s./(b1-s))
    input [N-1:0]b_xl ,          //параметр по входу x b - cередина сигмоиды
    input [N-1:0]b1_xl,          //параметр по входу x b1=s/(1-exp(-0.5))
    input [N-1:0]s_xl,            //параметр по входу x s - сигма сигмоиды 
    input [1:0]  ft_xl,          //тип активационной функции
	input [N-1:0]a0_yl,			//Коэффициент по входу y a0=sqrt(w_y)*sqrt(1-exp(-0.5))/s
	input [N-1:0]a1_yl,			//Коэффициент по входу y a1=sqrt(w_y)*sqrt((1-exp(-0.5))./s./(b1-s))
    input [N-1:0]b_yl ,          //параметр по входу y b - cередина сигмоиды
    input [N-1:0]b1_yl,          //параметр по входу y b1=s/(1-exp(-0.5))
    input [N-1:0]s_yl,            //параметр по входу x s - сигма сигмоиды 
    input [1:0]  ft_yl,          //тип активационной функции
    input [N-1:0]w_xl,           //весовой коэффициент по входу x [-1 1]
    input [N-1:0]w_yl,           //весовой коэффициент по входу y [-1 1]
//(правая функция принадлежноси) 
	input [N-1:0]a0_xr,			//Коэффициент по входу x a0=sqrt(w_x)*sqrt(1-exp(-0.5))/s
	input [N-1:0]a1_xr,			//Коэффициент по входу x a1=sqrt(w_x)*sqrt((1-exp(-0.5))./s./(b1-s))
    input [N-1:0]b_xr ,          //параметр по входу x b - cередина сигмоиды
    input [N-1:0]b1_xr,          //параметр по входу x b1=s/(1-exp(-0.5))
    input [N-1:0]s_xr,            //параметр по входу x s - сигма сигмоиды 
    input [1:0]  ft_xr,          //тип активационной функции
	input [N-1:0]a0_yr,			//Коэффициент по входу y a0=sqrt(w_y)*sqrt(1-exp(-0.5))/s
	input [N-1:0]a1_yr,			//Коэффициент по входу y a1=sqrt(w_y)*sqrt((1-exp(-0.5))./s./(b1-s))
    input [N-1:0]b_yr ,          //параметр по входу y b - cередина сигмоиды
    input [N-1:0]b1_yr,          //параметр по входу y b1=s/(1-exp(-0.5))
    input [N-1:0]s_yr,            //параметр по входу x s - сигма сигмоиды 
    input [1:0]  ft_yr,          //тип активационной функции
    input [N-1:0]w_xr,           //весовой коэффициент по входу x [-1 1]
    input [N-1:0]w_yr,           //весовой коэффициент по входу y [-1 1]
	output reg [N-1:0]out,          //Выход активационной функции
	output reg rdy			    	//Флаг окончания вычислений
	);


wire [N-1:0]ax_l;       //выход активационной функции входа x(левая функция принадлежности)
wire [N-1:0]ay_l;       //выход активационной функции входа y(левая функция принадлежности)
wire [N-1:0]ax_r;       //выход активационной функции входа x(правая функция принадлежности)
wire [N-1:0]ay_r;       //выход активационной функции входа y(правая функция принадлежности)
wire af_rdy;            //флаг готовности результата на выходе активационной функции


rbf_actfunc_cordic      //Активационная функция по входу x(левая функция принадлежности)
	#(.N(N), 			//Число бит входа и коэффициентов
      .bN(bN),           //Число бит целой части b,b1 и s  
      .aN(aN)
	) af_core_x_left
	(
	.rst(rst),			//Асинхронный сброс
	.clk(clk),			//Тактовый генератор
	.start(start),		//Строб старта
	.x(x),				//Вход [-1 1]
	.a0(a0_xl),			//Коэффициент a0=sqrt(w)*sqrt(1-exp(-0.5))/s
	.a1(a1_xl),			//Коэффициент a1=sqrt(w)*sqrt((1-exp(-0.5))./s./(b1-s))
    .b(b_xl),           //параметр b - середина сигмоиды
    .b1(b1_xl),         //параметр b1=s/(1-exp(-0.5))
    .s(s_xl),           //параметр s - сигма сигмоиды 
    .w(w_xl),           //весовой коэффициент [-1 1]
    .func_type(ft_xl),  //типа активационной функции    
	.y(ax_l),	 	    //Выход активационной функции в виде потока
	.rdy(af_rdy)	  	//Флаг выхода первого бита результата
	);

rbf_actfunc_cordic      //Активационная функция по входу x(правая функция принадлежности)
	#(.N(N), 			//Число бит входа и коэффициентов
      .bN(bN),          //Число бит целой части b,b1 и s  
      .aN(aN)
	) af_core_x_right
	(
	.rst(rst),			//Асинхронный сброс
	.clk(clk),			//Тактовый генератор
	.start(start),		//Строб старта
	.x(x),				//Вход [-1 1]
	.a0(a0_xr),			//Коэффициент a0=sqrt(w)*sqrt(1-exp(-0.5))/s
	.a1(a1_xr),			//Коэффициент a1=sqrt(w)*sqrt((1-exp(-0.5))./s./(b1-s))
    .b(b_xr),           //параметр b - середина сигмоиды
    .b1(b1_xr),         //параметр b1=s/(1-exp(-0.5))
    .s(s_xr),           //параметр s - сигма сигмоиды 
    .w(w_xr),           //весовой коэффициент [-1 1]
    .func_type(ft_xr),  //типа активационной функции    
  	.y(ax_r),	 	    //Выход активационной функции в виде потока
	.rdy()	  	//Флаг выхода первого бита результата
	);

rbf_actfunc_cordic      //Активационная функция по входу y(левая функция принадлежности)
	#(.N(N), 			//Число бит входа и коэффициентов
      .bN(bN),          //Число бит целой части b,b1 и s  
      .aN(aN)
	) af_core_y_left
	(
	.rst(rst),			//Асинхронный сброс
	.clk(clk),			//Тактовый генератор
	.start(start),		//Строб старта
	.x(y),				//Вход [-1 1]
	.a0(a0_yl),			//Коэффициент a0=sqrt(w)*sqrt(1-exp(-0.5))/s
	.a1(a1_yl),			//Коэффициент a1=sqrt(w)*sqrt((1-exp(-0.5))./s./(b1-s))
    .b(b_yl),           //параметр b - середина сигмоиды
    .b1(b1_yl),         //параметр b1=s/(1-exp(-0.5))
    .s(s_yl),           //параметр s - сигма сигмоиды 
    .w(w_yl),           //весовой коэффициент [-1 1]
    .func_type(ft_yl),  //типа активационной функции    
    
	.y(ay_l),	 	    //Выход активационной функции в виде потока
	.rdy()	  	//Флаг выхода первого бита результата
	);

rbf_actfunc_cordic      //Активационная функция по входу x(правая функция принадлежности)
	#(.N(N), 			//Число бит входа и коэффициентов
      .bN(bN),           //Число бит целой части b,b1 и s  
      .aN(aN)
	) af_core_y_right
	(
	.rst(rst),			//Асинхронный сброс
	.clk(clk),			//Тактовый генератор
	.start(start),		//Строб старта
	.x(y),				//Вход [-1 1]
	.a0(a0_yr),			//Коэффициент a0=sqrt(w)*sqrt(1-exp(-0.5))/s
	.a1(a1_yr),			//Коэффициент a1=sqrt(w)*sqrt((1-exp(-0.5))./s./(b1-s))
    .b(b_yr),           //параметр b - середина сигмоиды
    .b1(b1_yr),         //параметр b1=s/(1-exp(-0.5))
    .s(s_yr),           //параметр s - сигма сигмоиды 
    .w(w_yr),           //весовой коэффициент [-1 1]
    .func_type(ft_yr),  //типа активационной функции    
    
	.y(ay_r),	 	    //Выход активационной функции в виде потока
	.rdy()	  	//Флаг выхода первого бита результата
	);

reg start_c;   //Строб старта умножителя
reg [N-1:0]mult_a;  //множитель а
reg [N-1:0]mult_b;  //множитель b
wire [N-1:0]mult_c; //результат умножения
wire mult_rdy;       //флаг готовности результата


cordic_mult #(.N(N))                //Умножитель, реализующий правила
        fuzzy_multiplier
    (.clk(clk),
     .rst(rst),
     .a(mult_a),
     .b(mult_b),
     .start(start_c),
     .c(mult_c),
     .rdy(mult_rdy));

reg [N-1:0]y_left;  //результат перемножения левых термов по входу x и y

//typedef enum logic[2:0] {  
parameter
	st_idle			= 3'b001,
	st_mul_left		= 3'b010,
	st_mul_right	= 3'b100
	;//} MultState;
	
	reg [2:0] /*MultState*/ state;
always @(posedge clk, posedge rst)
    if(rst)
        begin
            mult_a <= 0;
            mult_b <= 0;
            start_c <= 0;
            state <=  st_idle;
            out <= 0;
            rdy <= 0;
            y_left <= 0;
        end else
        case (state)
            st_idle:
                begin
                    if(af_rdy)
                        begin   
                            mult_a<=ax_l;    //умножаем левые термы
                            mult_b<=ay_l;
                            start_c <= 1;
                            state <= st_mul_left;
                        end
                    rdy<=0;
                end
            st_mul_left:
                begin
                    if(mult_rdy)
                        begin
                            y_left <= mult_c;  //сохраняем результат умножения
                            mult_a<=ax_r;      //умножаем правые термы
                            mult_b<=ay_r;
                            start_c <= 1;
                            state <= st_mul_right;
                        end else
                            start_c <= 0;
                end
            st_mul_right:
                begin
                    if(mult_rdy)
                        begin
                            out <= mult_c - y_left;   //Выводим в результат разницу между правилами
                            rdy <=1;                  //выставляем флаг готовности
                            state <= st_idle;
                        end else
                            start_c <= 0;
                end
            
        endcase


endmodule

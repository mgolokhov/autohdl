`define test1 first_test
module inst1(
input a,
input b);
endmodule

module f2 ();

 f3 inst_f3();

endmodule
module f4_dsn1_tb();
endmodule
module inst2(
input a,
input b);
endmodule

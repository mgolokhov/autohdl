module f7();
endmodule

module f1_core2 ();
endmodule
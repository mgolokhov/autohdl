module non_top();
endmodule
module top(
input a,
output b
);

blk_mem_gen_v7_3 blk_mem_gen_v7_3_inst();


endmodule
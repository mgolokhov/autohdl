module f3_dsn1_uncopied();

endmodule
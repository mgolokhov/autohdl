module top_command_line();
endmodule
module f4();
f5 inst_f5();
f6 inst_f6();
//no inst_f7
endmodule

module f3 ();
f4 inst_f4();
endmodule